// Dataflow inverter
module not1_d (
  input  wire a,
  output wire y
);
  assign y = ~a;
endmodule

