// NOTE: This file is not used by the practice build.
// It remains here only as a scratchpad/open tab in your IDE.
// For interview-relevant modules and self-checking testbenches
// see the src/ and tb/ directories. If you want a 2:1 mux example,
// open src/dataflow/mux2_d.v or src/additions/gate/mux2_g.v.

/* Not used; keeping commented per your request
module mux2to1(
  input  wire a,
  input  wire b,
  input  wire sel,
  output wire y
);
  assign y = sel ? b : a;
endmodule
*/
