// Dataflow 2-input AND
module and2_d (
  input  wire a,
  input  wire b,
  output wire y
);
  assign y = a & b;
endmodule

